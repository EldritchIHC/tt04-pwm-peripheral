/*PWM Module 1*/
`define CONTROL_REG1 0
`define PERIOD_MSB1 1
`define PERIOD_LSB1 2
`define ACTION_REG_A1 3
`define COMP_A_MSB_A1 4
`define COMP_A_LSB_A1 5
`define COMP_A_MSB_B1 6
`define COMP_A_LSB_B1 7
`define DEADBAND_REG_A1 8
`define ACTION_REG_B1 9
`define COMP_B_MSB_A1 10
`define COMP_B_LSB_A1 11
`define COMP_B_MSB_B1 12
`define COMP_B_LSB_B1 13
`define DEADBAND_REG_B1 14
/*PWM Module 2*/
`define CONTROL_REG2 15
`define PERIOD_MSB2 16
`define PERIOD_LSB2 17
`define PHASE_MSB2  18
`define PHASE_LSB2  19
`define ACTION_REG_A2 20
`define COMP_A_MSB_A2 21
`define COMP_A_LSB_A2 22
`define COMP_A_MSB_B2 23
`define COMP_A_LSB_B2 24
`define DEADBAND_REG_A2 25
`define ACTION_REG_B2 26
`define COMP_B_MSB_A2 27
`define COMP_B_LSB_A2 28
`define COMP_B_MSB_B2 29
`define COMP_B_LSB_B2 30
`define DEADBAND_REG_B2 31
/*PWM Module 3*/
`define CONTROL_REG3 32
`define PERIOD_MSB3 33
`define PERIOD_LSB3 34
`define PHASE_MSB3  35
`define PHASE_LSB3  36
`define ACTION_REG_A3 37
`define COMP_A_MSB_A3 38
`define COMP_A_LSB_A3 39
`define COMP_A_MSB_B3 40
`define COMP_A_LSB_B3 41
`define DEADBAND_REG_A3 42
`define ACTION_REG_B3 43
`define COMP_B_MSB_A3 44
`define COMP_B_LSB_A3 45
`define COMP_B_MSB_B3 46
`define COMP_B_LSB_B3 47
`define DEADBAND_REG_B3 48